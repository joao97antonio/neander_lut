library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use ieee.std_logic_unsigned.all;
use ieee.std_logic_arith.all;
use IEEE.STD_LOGIC_1164.ALL;

entity lut_sub is
    port(
        input_lut : in std_logic_vector(7 downto 0);
        output_lut : in std_logic_vector(3 downto 0)
    );
end lut_mult;
architecture behavior of lut_sub is
        
        type lut is array (integer range 0 to 255) of std_logic_vector(3 downto 0); 
        signal sub_lut : lut;
        signal output_4bits : in std_logic_vector(7 downto 0);
        
        begin
        output_4bits <= add_lut(conv_integer(input_lut));
        
        mult_lut (0)<= "00000000";
		mult_lut (1)<= "00000000";
		mult_lut (2)<= "00000000";
		mult_lut (3)<= "00000000";
		mult_lut (4)<= "00000000";
		mult_lut (5)<= "00000000";
		mult_lut (6)<= "00000000";
		mult_lut (7)<= "00000000";
   	    mult_lut (8)<= "00000000";
		mult_lut (9)<= "00000000";
		mult_lut (10)<= "00000000";
		mult_lut (11)<= "00000000";
		mult_lut (12)<= "00000000";
		mult_lut (13)<= "00000000";
		mult_lut (14)<= "00000000";
		mult_lut (15)<= "00000000";
        mult_lut (16)<= "00000000";
		mult_lut (17)<= "00000001";
		mult_lut (18)<= "00000010";
		mult_lut (19)<= "00000011";
		mult_lut (20)<= "00000100";
		mult_lut (21)<= "00000101";
		mult_lut (22)<= "00000110";
		mult_lut (23)<= "00000111";
   	    mult_lut (24)<= "00001000";
		mult_lut (25)<= "00001001";
		mult_lut (26)<= "00001010";
		mult_lut (27)<= "00001011";
		mult_lut (28)<= "00001100";
		mult_lut (29)<= "00001101";
		mult_lut (30)<= "00001110";
		mult_lut (31)<= "00001111";
        mult_lut (32)<= "00000000";
		mult_lut (33)<= "00000010";
		mult_lut (34)<= "00000100";
		mult_lut (35)<= "00000110";
		mult_lut (36)<= "00001000";
		mult_lut (37)<= "00001010";
		mult_lut (38)<= "00001100";
		mult_lut (39)<= "00001110";
   	    mult_lut (40)<= "00010000";
		mult_lut (41)<= "00010010";
		mult_lut (42)<= "00010100";
		mult_lut (43)<= "00010110";
		mult_lut (44)<= "00011000";
		mult_lut (45)<= "00011010";
		mult_lut (46)<= "00011100";
		mult_lut (47)<= "00011110";
        mult_lut (48)<= "00000000";
		mult_lut (49)<= "00000011";
		mult_lut (50)<= "00000110";
		mult_lut (51)<= "00001001";
		mult_lut (52)<= "00001100";
		mult_lut (53)<= "00001111";
		mult_lut (54)<= "00010010";
		mult_lut (55)<= "00010101";
   	    mult_lut (56)<= "00011000";
		mult_lut (57)<= "00011011";
		mult_lut (58)<= "00011110";
		mult_lut (59)<= "00100001";
		mult_lut (60)<= "00100100";
		mult_lut (61)<= "00100111";
		mult_lut (62)<= "00101010";
		mult_lut (63)<= "00101101";
        mult_lut (64)<= "00000000";
		mult_lut (65)<= "00000100";
		mult_lut (66)<= "00001000";
		mult_lut (67)<= "00001100";
		mult_lut (68)<= "00010000";
		mult_lut (69)<= "00010100";
		mult_lut (70)<= "00011000";
		mult_lut (71)<= "00011100";
   	    mult_lut (72)<= "00100000";
		mult_lut (73)<= "00100100";
		mult_lut (74)<= "00101000";
		mult_lut (75)<= "00101100";
		mult_lut (76)<= "00110000";
		mult_lut (77)<= "00110100";
		mult_lut (78)<= "00111000";
		mult_lut (79)<= "00111100";
        mult_lut (80)<= "00000000";
		mult_lut (81)<= "00000101";
		mult_lut (82)<= "00001010";
		mult_lut (83)<= "00001111";
		mult_lut (84)<= "00010100";
		mult_lut (85)<= "00011001";
		mult_lut (86)<= "00011110";
		mult_lut (87)<= "00100011";
   	    mult_lut (88)<= "00101000";
		mult_lut (89)<= "00101101";
		mult_lut (90)<= "00110010";
		mult_lut (91)<= "00110111";
		mult_lut (92)<= "00111100";
		mult_lut (93)<= "01000001";
		mult_lut (94)<= "01000110";
		mult_lut (95)<= "01001011";
        mult_lut (96)<= "00000000";
		mult_lut (97)<= "00000110";
		mult_lut (98)<= "00001100";
		mult_lut (99)<= "00010010";
		mult_lut (100)<= "00011000";
		mult_lut (101)<= "00011110";
		mult_lut (102)<= "00100100";
		mult_lut (103)<= "00101010";
   	    mult_lut (104)<= "00110000";
		mult_lut (105)<= "00110110";
		mult_lut (106)<= "00111100";
		mult_lut (107)<= "01000010";
		mult_lut (108)<= "01001000";
		mult_lut (109)<= "01001110";
		mult_lut (110)<= "01010100";
		mult_lut (111)<= "01011010";
        mult_lut (112)<= "00000000";
		mult_lut (113)<= "00000111";
		mult_lut (114)<= "00001110";
		mult_lut (115)<= "00010101";
		mult_lut (116)<= "00011100";
		mult_lut (117)<= "00100011";
		mult_lut (118)<= "00101010";
		mult_lut (119)<= "00110001";
   	    mult_lut (120)<= "00111000";
		mult_lut (121)<= "00111111";
		mult_lut (122)<= "01000110";
		mult_lut (123)<= "01001101";
		mult_lut (124)<= "01010100";
		mult_lut (125)<= "01011011";
		mult_lut (126)<= "01100010";
		mult_lut (127)<= "01101001";
        mult_lut (128)<= "00000000";
		mult_lut (129)<= "00001000";
		mult_lut (130)<= "00010000";
		mult_lut (131)<= "00011000";
		mult_lut (132)<= "00100000";
		mult_lut (133)<= "00101000";
		mult_lut (134)<= "00110000";
		mult_lut (135)<= "00111000";
   	    mult_lut (136)<= "01000000";
		mult_lut (137)<= "01001000";
		mult_lut (138)<= "01010000";
		mult_lut (139)<= "01011000";
		mult_lut (140)<= "01100000";
		mult_lut (141)<= "01101000";
		mult_lut (142)<= "01110000";
		mult_lut (143)<= "01111000";
        mult_lut (144)<= "00000000";
		mult_lut (145)<= "00001001";
		mult_lut (146)<= "00010010";
		mult_lut (147)<= "00011011";
		mult_lut (148)<= "00100100";
		mult_lut (149)<= "00101101";
		mult_lut (150)<= "00110110";
		mult_lut (151)<= "00111111";
   	    mult_lut (152)<= "01001000";
		mult_lut (153)<= "01010001";
		mult_lut (154)<= "01011010";
		mult_lut (155)<= "01100011";
		mult_lut (156)<= "01101100";
		mult_lut (157)<= "01110101";
		mult_lut (158)<= "01111110";
		mult_lut (159)<= "10000111";
        mult_lut (160)<= "00000000";
		mult_lut (161)<= "00001010";
		mult_lut (162)<= "00010100";
		mult_lut (163)<= "00011110";
		mult_lut (164)<= "00101000";
		mult_lut (165)<= "00110010";
		mult_lut (166)<= "00111100";
		mult_lut (167)<= "01000110";
   	    mult_lut (168)<= "01010000";
		mult_lut (169)<= "01011010";
		mult_lut (170)<= "01100100";
		mult_lut (171)<= "01101110";
		mult_lut (172)<= "01111000";
		mult_lut (173)<= "10000010";
		mult_lut (174)<= "10001100";
		mult_lut (175)<= "10010110";
        mult_lut (176)<= "00000000";
		mult_lut (177)<= "00001011";
		mult_lut (178)<= "00010110";
		mult_lut (179)<= "00100001";
		mult_lut (180)<= "00101100";
		mult_lut (181)<= "00110111";
		mult_lut (182)<= "01000010";
		mult_lut (183)<= "01001101";
   	    mult_lut (184)<= "01011000";
		mult_lut (185)<= "01100011";
		mult_lut (186)<= "01101110";
		mult_lut (187)<= "01111001";
		mult_lut (188)<= "10000100";
		mult_lut (189)<= "10001111";
		mult_lut (190)<= "10011010";
		mult_lut (191)<= "10100101";
        mult_lut (192)<= "00000000";
		mult_lut (193)<= "00001100";
		mult_lut (194)<= "00011000";
		mult_lut (195)<= "00100100";
		mult_lut (196)<= "00110000";
		mult_lut (197)<= "00111100";
		mult_lut (198)<= "01001000";
		mult_lut (199)<= "01010100";
   	    mult_lut (200)<= "01100000";
		mult_lut (201)<= "01101100";
		mult_lut (202)<= "01111000";
		mult_lut (203)<= "10000100";
		mult_lut (204)<= "10010000";
		mult_lut (205)<= "10011100";
		mult_lut (206)<= "10101000";
		mult_lut (207)<= "10110100";
        mult_lut (208)<= "00000000";
		mult_lut (209)<= "00001101";
		mult_lut (210)<= "00011010";
		mult_lut (211)<= "00100111";
		mult_lut (212)<= "00110100";
		mult_lut (213)<= "01000001";
		mult_lut (214)<= "01001110";
		mult_lut (215)<= "01011011";
   	    mult_lut (216)<= "01101000";
		mult_lut (217)<= "01110101";
		mult_lut (218)<= "10000010";
		mult_lut (219)<= "10001111";
		mult_lut (220)<= "10011100";
		mult_lut (221)<= "10101001";
		mult_lut (222)<= "10110110";
		mult_lut (223)<= "11000011";
        mult_lut (224)<= "00000000";
		mult_lut (225)<= "00001110";
		mult_lut (226)<= "00011100";
		mult_lut (227)<= "00101010";
		mult_lut (228)<= "00111000";
		mult_lut (229)<= "01000110";
		mult_lut (230)<= "01010100";
		mult_lut (231)<= "01100010";
   	    mult_lut (232)<= "01110000";
		mult_lut (233)<= "01111110";
		mult_lut (234)<= "10001100";
		mult_lut (235)<= "10011010";
		mult_lut (236)<= "10101000";
		mult_lut (237)<= "10110110";
		mult_lut (238)<= "11000100";
		mult_lut (239)<= "11010010";
        mult_lut (240)<= "00000000";
		mult_lut (241)<= "00001111";
		mult_lut (242)<= "00011110";
		mult_lut (243)<= "00101101";
		mult_lut (244)<= "00111100";
		mult_lut (245)<= "01001011";
		mult_lut (246)<= "01011010";
		mult_lut (247)<= "01101001";
   	    mult_lut (248)<= "01111000";
		mult_lut (249)<= "10000111";
		mult_lut (250)<= "10010110";
		mult_lut (251)<= "10100101";
		mult_lut (252)<= "10110100";
		mult_lut (253)<= "11000011";
		mult_lut (254)<= "11010010";
		mult_lut (255)<= "11100001"; 

    output_lut <= output_4bits(3 downto 0);
end behavior;